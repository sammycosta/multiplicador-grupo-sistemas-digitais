library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity somador is
    generic(N: integer);
	port(A, B: in std_logic_vector(N-1 downto 0);
		S: out std_logic_vector(N-1 downto 0));
end somador;

architecture arch of somador is
    -- somador comportamental
begin
    S <= A + B;
end arch;
